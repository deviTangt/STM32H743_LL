//********************************//
//! ģ��: spi_test
//  ����: spi_master��spi_slave����ģ��
//********************************//
module spi_test(
    input  wire                     sys_clk         ,   //? ϵͳʱ��
    input  wire                     sys_rst_n       ,   //? ϵͳ��λ������Ч

    input  wire                     en_spi    
);

//**************************************// ������д         //**********************************//


//**************************************// �ź�����         //**********************************//
wire                cs;
wire                sclk;
wire                mosi;
wire                miso;

wire                wr_ack;
wire                re_ack;

wire    [7 : 0]     master_rx;
wire    [7 : 0]     slave_rx;

wire                cs_ctrl;
assign              cs_ctrl = en_spi;

//**************************************// �������         //**********************************//



//**************************************// ��ģ�����       //**********************************//
spi_master#(
	.CPOL           (1'b1)					    ,			// ʱ�Ӽ��Կ���
	.CPHA           (1'b1)									// ʱ����λ����
)
ins_spi_master
(	
	.sys_clk		(sys_clk)                   ,     	    // ʱ���ź�
	.sys_rst_n		(sys_rst_n)                 ,   		// ��λ�ź�

	.cs				(cs)                        ,           // Ƭѡ�ź�
	.sclk			(sclk)                      ,        	// ʱ���ź����
	.mosi			(mosi)                      ,        	// ���豸������豸����������
	.miso			(miso)                      ,        	// ���豸������豸���������

	.cs_ctrl		(cs_ctrl)                   ,     	    // Ƭѡ�����ź� cs = cs_ctrl
	.clk_div_val	(50 - 1)                    ,           // ʱ�ӷ�Ƶֵ 1M

	.wr_req			(en_spi)                    ,      	    // д�����ź�
	.wr_ack			(wr_ack)                    ,      	    // дӦ���ź�

	.data_tx		(master_rx + 8'b1)          ,           // ��������
	.data_rx 		(master_rx)                             // �������
);

spi_slave#(
	.CPOL           (1'b1)					    ,			// ʱ�Ӽ��Կ���
	.CPHA           (1'b1)								    // ʱ����λ����
)
ins_spi_slave
(	
	.sys_clk		(sys_clk)                   ,     	    // ʱ���ź�
	.sys_rst_n		(sys_rst_n)                 ,   	    // ��λ�ź�
                           
	.cs				(cs)                        ,           // Ƭѡ�ź�
	.sclk			(sclk)                      ,           // ʱ���ź����
	.mosi			(mosi)                      ,           // ���豸������豸����������
	.miso			(miso)                      ,           // ���豸������豸���������
                            
	.re_ack			(re_ack)                    ,      	    // ��Ӧ���ź�
                             
	.data_tx		(slave_rx + 8'd2)           ,           // ��������
	.data_rx 		(slave_rx)                              // �������
);  
//**************************************// ģ�����         //**********************************//
endmodule
