//********************************//
//! ģ��: spi_test
//  ����: spi_master��spi_slave����ģ��
//********************************//
module spi_test(
    input  wire                     sys_clk         ,   //? ϵͳʱ��
    input  wire                     sys_rst_n           //? ϵͳ��λ������Ч
);

//**************************************// ������д         //**********************************//


//**************************************// �ź�����         //**********************************//
wire                cs;
wire                sclk;
wire                mosi;
wire                miso;

//**************************************// �������         //**********************************//



//**************************************// ��ģ�����       //**********************************//
spi_master#(
	.CPOL           (1'b1)						,			// ʱ�Ӽ��Կ���
	.CPHA           (1'b1)									// ʱ����λ����
)
ins_spi_master
(	
	.sys_clk		(sys_clk)                          ,     		// ʱ���ź�
	.sys_rst_n		(sys_rst_n)                          ,   		// ��λ�ź�
                    
	.cs				(cs)                          ,          	// Ƭѡ�ź�
	.sclk			(sclk)                          ,        	// ʱ���ź����
	.mosi			(mosi)                          ,        	// ���豸������豸����������
	.miso			(miso)                          ,        	// ���豸������豸���������
                         
	.cs_ctrl		()                          ,     		// Ƭѡ�����ź� cs = cs_ctrl
	.clk_div_val	()                          ,          	// ʱ�ӷ�Ƶֵ
                     
	.wr_req			()                          ,      		// д�����ź�
	.wr_ack			()                          ,      		// дӦ���ź�
                      
	.data_tx		()                          ,           // ��������
	.data_rx 		()                                     	// �������
);

spi_slave#(
	.CPOL               (1'b1)					,			// ʱ�Ӽ��Կ���
	.CPHA               (1'b1)								// ʱ����λ����
)
ins_spi_slave
(	
	.sys_clk		(sys_clk)                          ,     	    // ʱ���ź�
	.sys_rst_n		(sys_rst_n)                          ,   	    // ��λ�ź�
                           
	.cs				(cs)                          ,           // Ƭѡ�ź�
	.sclk			(sclk)                          ,           // ʱ���ź����
	.mosi			(mosi)                          ,           // ���豸������豸����������
	.miso			(miso)                          ,           // ���豸������豸���������
                    
	.clk_div_val	()                          ,           // ʱ�ӷ�Ƶֵ
                            
	.re_ack			()                          ,      	    // ��Ӧ���ź�
                             
	.data_tx		()                          ,           // ��������
	.data_rx 		()                                      // �������
);  
//**************************************// ģ�����         //**********************************//
endmodule
